`timescale 1ns/1ns

module alu_tb;
	reg [11:0]x;
	reg [11:0]y;
    reg [2:0]op;
	wire [11:0]z;
	alu u1 (.op(op), .op1(x), .op2(y), .out(z));
	initial begin
		$dumpfile("alu_tb.vcd");
		$dumpvars(0, alu_tb);
        $monitor("X=%b, Y=%b, OP=%b, Z=%b", x, y, op, z);
		x=12'b001111100000; y=12'b001111100000; op=3'b000; #20;
		x=12'b000000001111; y=12'b000000000011; op=3'b001; #20;
		x=12'b000000001111; y=12'b000000000011; op=3'b010; #20;
		x=12'b000000001111; y=12'b000000000011; op=3'b011; #20;
		x=12'b000000001111; y=12'b000000000011; op=3'b100; #20;
		x=12'b010000100000; y=12'b001111000000; op=3'b101; #20;
		x=12'b010000100000; y=12'b001111000000; op=3'b110; #20;
		x=12'b000000001111; y=12'b000000001111; op=3'b111; #20;
	end
	
endmodule
